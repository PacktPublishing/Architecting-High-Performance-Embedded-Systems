-- Load the standard libraries

library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;

-- Define the 4-bit adder inputs and outputs

entity ADDER4LUT is
  port (
    A4     : in    std_logic_vector(3 downto 0);
    B4     : in    std_logic_vector(3 downto 0);
    SUM4   : out   std_logic_vector(3 downto 0);
    C_OUT4 : out   std_logic
  );
end entity ADDER4LUT;

-- Define the behavior of the 4-bit adder

architecture BEHAVIORAL of ADDER4LUT is

begin

  ADDER_LUT : process (A4, B4) is

    variable concat_input : std_logic_vector(7 downto 0);

  begin

    concat_input := A4 & B4;

    case concat_input is

      when "00000000" =>
        SUM4 <= "0000"; C_OUT4 <= '0';
      when "00000001" =>
        SUM4 <= "0001"; C_OUT4 <= '0';
      when "00000010" =>
        SUM4 <= "0010"; C_OUT4 <= '0';
      when "00000011" =>
        SUM4 <= "0011"; C_OUT4 <= '0';
      when "00000100" =>
        SUM4 <= "0100"; C_OUT4 <= '0';
      when "00000101" =>
        SUM4 <= "0101"; C_OUT4 <= '0';
      when "00000110" =>
        SUM4 <= "0110"; C_OUT4 <= '0';
      when "00000111" =>
        SUM4 <= "0111"; C_OUT4 <= '0';
      when "00001000" =>
        SUM4 <= "1000"; C_OUT4 <= '0';
      when "00001001" =>
        SUM4 <= "1001"; C_OUT4 <= '0';
      when "00001010" =>
        SUM4 <= "1010"; C_OUT4 <= '0';
      when "00001011" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "00001100" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "00001101" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "00001110" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "00001111" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "00010000" =>
        SUM4 <= "0001"; C_OUT4 <= '0';
      when "00010001" =>
        SUM4 <= "0010"; C_OUT4 <= '0';
      when "00010010" =>
        SUM4 <= "0011"; C_OUT4 <= '0';
      when "00010011" =>
        SUM4 <= "0100"; C_OUT4 <= '0';
      when "00010100" =>
        SUM4 <= "0101"; C_OUT4 <= '0';
      when "00010101" =>
        SUM4 <= "0110"; C_OUT4 <= '0';
      when "00010110" =>
        SUM4 <= "0111"; C_OUT4 <= '0';
      when "00010111" =>
        SUM4 <= "1000"; C_OUT4 <= '0';
      when "00011000" =>
        SUM4 <= "1001"; C_OUT4 <= '0';
      when "00011001" =>
        SUM4 <= "1010"; C_OUT4 <= '0';
      when "00011010" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "00011011" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "00011100" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "00011101" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "00011110" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "00011111" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "00100000" =>
        SUM4 <= "0010"; C_OUT4 <= '0';
      when "00100001" =>
        SUM4 <= "0011"; C_OUT4 <= '0';
      when "00100010" =>
        SUM4 <= "0100"; C_OUT4 <= '0';
      when "00100011" =>
        SUM4 <= "0101"; C_OUT4 <= '0';
      when "00100100" =>
        SUM4 <= "0110"; C_OUT4 <= '0';
      when "00100101" =>
        SUM4 <= "0111"; C_OUT4 <= '0';
      when "00100110" =>
        SUM4 <= "1000"; C_OUT4 <= '0';
      when "00100111" =>
        SUM4 <= "1001"; C_OUT4 <= '0';
      when "00101000" =>
        SUM4 <= "1010"; C_OUT4 <= '0';
      when "00101001" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "00101010" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "00101011" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "00101100" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "00101101" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "00101110" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "00101111" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "00110000" =>
        SUM4 <= "0011"; C_OUT4 <= '0';
      when "00110001" =>
        SUM4 <= "0100"; C_OUT4 <= '0';
      when "00110010" =>
        SUM4 <= "0101"; C_OUT4 <= '0';
      when "00110011" =>
        SUM4 <= "0110"; C_OUT4 <= '0';
      when "00110100" =>
        SUM4 <= "0111"; C_OUT4 <= '0';
      when "00110101" =>
        SUM4 <= "1000"; C_OUT4 <= '0';
      when "00110110" =>
        SUM4 <= "1001"; C_OUT4 <= '0';
      when "00110111" =>
        SUM4 <= "1010"; C_OUT4 <= '0';
      when "00111000" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "00111001" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "00111010" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "00111011" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "00111100" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "00111101" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "00111110" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "00111111" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "01000000" =>
        SUM4 <= "0100"; C_OUT4 <= '0';
      when "01000001" =>
        SUM4 <= "0101"; C_OUT4 <= '0';
      when "01000010" =>
        SUM4 <= "0110"; C_OUT4 <= '0';
      when "01000011" =>
        SUM4 <= "0111"; C_OUT4 <= '0';
      when "01000100" =>
        SUM4 <= "1000"; C_OUT4 <= '0';
      when "01000101" =>
        SUM4 <= "1001"; C_OUT4 <= '0';
      when "01000110" =>
        SUM4 <= "1010"; C_OUT4 <= '0';
      when "01000111" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "01001000" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "01001001" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "01001010" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "01001011" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "01001100" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "01001101" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "01001110" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "01001111" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "01010000" =>
        SUM4 <= "0101"; C_OUT4 <= '0';
      when "01010001" =>
        SUM4 <= "0110"; C_OUT4 <= '0';
      when "01010010" =>
        SUM4 <= "0111"; C_OUT4 <= '0';
      when "01010011" =>
        SUM4 <= "1000"; C_OUT4 <= '0';
      when "01010100" =>
        SUM4 <= "1001"; C_OUT4 <= '0';
      when "01010101" =>
        SUM4 <= "1010"; C_OUT4 <= '0';
      when "01010110" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "01010111" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "01011000" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "01011001" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "01011010" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "01011011" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "01011100" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "01011101" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "01011110" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "01011111" =>
        SUM4 <= "0100"; C_OUT4 <= '1';
      when "01100000" =>
        SUM4 <= "0110"; C_OUT4 <= '0';
      when "01100001" =>
        SUM4 <= "0111"; C_OUT4 <= '0';
      when "01100010" =>
        SUM4 <= "1000"; C_OUT4 <= '0';
      when "01100011" =>
        SUM4 <= "1001"; C_OUT4 <= '0';
      when "01100100" =>
        SUM4 <= "1010"; C_OUT4 <= '0';
      when "01100101" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "01100110" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "01100111" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "01101000" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "01101001" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "01101010" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "01101011" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "01101100" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "01101101" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "01101110" =>
        SUM4 <= "0100"; C_OUT4 <= '1';
      when "01101111" =>
        SUM4 <= "0101"; C_OUT4 <= '1';
      when "01110000" =>
        SUM4 <= "0111"; C_OUT4 <= '0';
      when "01110001" =>
        SUM4 <= "1000"; C_OUT4 <= '0';
      when "01110010" =>
        SUM4 <= "1001"; C_OUT4 <= '0';
      when "01110011" =>
        SUM4 <= "1010"; C_OUT4 <= '0';
      when "01110100" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "01110101" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "01110110" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "01110111" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "01111000" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "01111001" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "01111010" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "01111011" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "01111100" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "01111101" =>
        SUM4 <= "0100"; C_OUT4 <= '1';
      when "01111110" =>
        SUM4 <= "0101"; C_OUT4 <= '1';
      when "01111111" =>
        SUM4 <= "0110"; C_OUT4 <= '1';
      when "10000000" =>
        SUM4 <= "1000"; C_OUT4 <= '0';
      when "10000001" =>
        SUM4 <= "1001"; C_OUT4 <= '0';
      when "10000010" =>
        SUM4 <= "1010"; C_OUT4 <= '0';
      when "10000011" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "10000100" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "10000101" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "10000110" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "10000111" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "10001000" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "10001001" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "10001010" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "10001011" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "10001100" =>
        SUM4 <= "0100"; C_OUT4 <= '1';
      when "10001101" =>
        SUM4 <= "0101"; C_OUT4 <= '1';
      when "10001110" =>
        SUM4 <= "0110"; C_OUT4 <= '1';
      when "10001111" =>
        SUM4 <= "0111"; C_OUT4 <= '1';
      when "10010000" =>
        SUM4 <= "1001"; C_OUT4 <= '0';
      when "10010001" =>
        SUM4 <= "1010"; C_OUT4 <= '0';
      when "10010010" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "10010011" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "10010100" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "10010101" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "10010110" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "10010111" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "10011000" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "10011001" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "10011010" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "10011011" =>
        SUM4 <= "0100"; C_OUT4 <= '1';
      when "10011100" =>
        SUM4 <= "0101"; C_OUT4 <= '1';
      when "10011101" =>
        SUM4 <= "0110"; C_OUT4 <= '1';
      when "10011110" =>
        SUM4 <= "0111"; C_OUT4 <= '1';
      when "10011111" =>
        SUM4 <= "1000"; C_OUT4 <= '1';
      when "10100000" =>
        SUM4 <= "1010"; C_OUT4 <= '0';
      when "10100001" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "10100010" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "10100011" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "10100100" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "10100101" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "10100110" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "10100111" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "10101000" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "10101001" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "10101010" =>
        SUM4 <= "0100"; C_OUT4 <= '1';
      when "10101011" =>
        SUM4 <= "0101"; C_OUT4 <= '1';
      when "10101100" =>
        SUM4 <= "0110"; C_OUT4 <= '1';
      when "10101101" =>
        SUM4 <= "0111"; C_OUT4 <= '1';
      when "10101110" =>
        SUM4 <= "1000"; C_OUT4 <= '1';
      when "10101111" =>
        SUM4 <= "1001"; C_OUT4 <= '1';
      when "10110000" =>
        SUM4 <= "1011"; C_OUT4 <= '0';
      when "10110001" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "10110010" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "10110011" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "10110100" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "10110101" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "10110110" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "10110111" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "10111000" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "10111001" =>
        SUM4 <= "0100"; C_OUT4 <= '1';
      when "10111010" =>
        SUM4 <= "0101"; C_OUT4 <= '1';
      when "10111011" =>
        SUM4 <= "0110"; C_OUT4 <= '1';
      when "10111100" =>
        SUM4 <= "0111"; C_OUT4 <= '1';
      when "10111101" =>
        SUM4 <= "1000"; C_OUT4 <= '1';
      when "10111110" =>
        SUM4 <= "1001"; C_OUT4 <= '1';
      when "10111111" =>
        SUM4 <= "1010"; C_OUT4 <= '1';
      when "11000000" =>
        SUM4 <= "1100"; C_OUT4 <= '0';
      when "11000001" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "11000010" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "11000011" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "11000100" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "11000101" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "11000110" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "11000111" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "11001000" =>
        SUM4 <= "0100"; C_OUT4 <= '1';
      when "11001001" =>
        SUM4 <= "0101"; C_OUT4 <= '1';
      when "11001010" =>
        SUM4 <= "0110"; C_OUT4 <= '1';
      when "11001011" =>
        SUM4 <= "0111"; C_OUT4 <= '1';
      when "11001100" =>
        SUM4 <= "1000"; C_OUT4 <= '1';
      when "11001101" =>
        SUM4 <= "1001"; C_OUT4 <= '1';
      when "11001110" =>
        SUM4 <= "1010"; C_OUT4 <= '1';
      when "11001111" =>
        SUM4 <= "1011"; C_OUT4 <= '1';
      when "11010000" =>
        SUM4 <= "1101"; C_OUT4 <= '0';
      when "11010001" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "11010010" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "11010011" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "11010100" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "11010101" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "11010110" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "11010111" =>
        SUM4 <= "0100"; C_OUT4 <= '1';
      when "11011000" =>
        SUM4 <= "0101"; C_OUT4 <= '1';
      when "11011001" =>
        SUM4 <= "0110"; C_OUT4 <= '1';
      when "11011010" =>
        SUM4 <= "0111"; C_OUT4 <= '1';
      when "11011011" =>
        SUM4 <= "1000"; C_OUT4 <= '1';
      when "11011100" =>
        SUM4 <= "1001"; C_OUT4 <= '1';
      when "11011101" =>
        SUM4 <= "1010"; C_OUT4 <= '1';
      when "11011110" =>
        SUM4 <= "1011"; C_OUT4 <= '1';
      when "11011111" =>
        SUM4 <= "1100"; C_OUT4 <= '1';
      when "11100000" =>
        SUM4 <= "1110"; C_OUT4 <= '0';
      when "11100001" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "11100010" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "11100011" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "11100100" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "11100101" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "11100110" =>
        SUM4 <= "0100"; C_OUT4 <= '1';
      when "11100111" =>
        SUM4 <= "0101"; C_OUT4 <= '1';
      when "11101000" =>
        SUM4 <= "0110"; C_OUT4 <= '1';
      when "11101001" =>
        SUM4 <= "0111"; C_OUT4 <= '1';
      when "11101010" =>
        SUM4 <= "1000"; C_OUT4 <= '1';
      when "11101011" =>
        SUM4 <= "1001"; C_OUT4 <= '1';
      when "11101100" =>
        SUM4 <= "1010"; C_OUT4 <= '1';
      when "11101101" =>
        SUM4 <= "1011"; C_OUT4 <= '1';
      when "11101110" =>
        SUM4 <= "1100"; C_OUT4 <= '1';
      when "11101111" =>
        SUM4 <= "1101"; C_OUT4 <= '1';
      when "11110000" =>
        SUM4 <= "1111"; C_OUT4 <= '0';
      when "11110001" =>
        SUM4 <= "0000"; C_OUT4 <= '1';
      when "11110010" =>
        SUM4 <= "0001"; C_OUT4 <= '1';
      when "11110011" =>
        SUM4 <= "0010"; C_OUT4 <= '1';
      when "11110100" =>
        SUM4 <= "0011"; C_OUT4 <= '1';
      when "11110101" =>
        SUM4 <= "0100"; C_OUT4 <= '1';
      when "11110110" =>
        SUM4 <= "0101"; C_OUT4 <= '1';
      when "11110111" =>
        SUM4 <= "0110"; C_OUT4 <= '1';
      when "11111000" =>
        SUM4 <= "0111"; C_OUT4 <= '1';
      when "11111001" =>
        SUM4 <= "1000"; C_OUT4 <= '1';
      when "11111010" =>
        SUM4 <= "1001"; C_OUT4 <= '1';
      when "11111011" =>
        SUM4 <= "1010"; C_OUT4 <= '1';
      when "11111100" =>
        SUM4 <= "1011"; C_OUT4 <= '1';
      when "11111101" =>
        SUM4 <= "1100"; C_OUT4 <= '1';
      when "11111110" =>
        SUM4 <= "1101"; C_OUT4 <= '1';
      when "11111111" =>
        SUM4 <= "1110"; C_OUT4 <= '1';
      when others =>
        SUM4 <= "UUUU"; C_OUT4 <= 'U';

    end case;

  end process ADDER_LUT;

end architecture BEHAVIORAL;
